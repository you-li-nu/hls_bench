
package vvectors is 
  subtype bit32 is integer;
  subtype bit4 is integer range 0 to 15;
  subtype bit16 is integer range 0 to 65535;
end vvectors;

